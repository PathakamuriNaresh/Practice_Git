hello all welcome to git lesson for practice to understand the basics of it
so here also in erh.sv the file is edited from the git
