hello everyone good to see you again
