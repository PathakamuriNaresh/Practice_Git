this file is added for the new branch1
