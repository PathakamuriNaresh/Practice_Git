hello all welcome to git lesson for practice
