new file added here
this new file is edited from the git 
