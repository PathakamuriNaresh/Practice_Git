hello all welcome to git lesson for practice to understand the basics of it
